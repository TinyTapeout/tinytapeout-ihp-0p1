`default_nettype none

module tt_logo ();
endmodule
